module Condition_Check (
    input [3:0] Cond, status,
    output is_valid
);
    
endmodule