module IF_Stage (
    input clk, rst, freeze, Branch_taken,
    input[31:0] BranchAddr,
    output reg [31:0] PC, 
	output[31:0] Instruction
);

wire[31:0] mem[0:46];
assign mem[0] = 32'b11100011101000000000000000010100; //MOV R0 ,#20 //R0 = 20
assign mem[1] = 32'b11100011101000000001101000000001; //MOV R1 ,#4096 //R1 = 4096
assign mem[2] = 32'b11100011101000000010000100000011; //MOV R2 ,#0xC0000000 //R2 = -1073741824
assign mem[3] = 32'b11100000100100100011000000000010; //ADDS R3 ,R2,R2 //R3 = -2147483648 
assign mem[4] = 32'b11100000101000000100000000000000; //ADC R4 ,R0,R0 //R4 = 41
assign mem[5] = 32'b11100000010001000101000100000100; //SUB R5 ,R4,R4,LSL #2 //R5 = -123
assign mem[6] = 32'b11100000110000000110000010100000; //SBC R6 ,R0,R0,LSR #1 //R6 = 10
assign mem[7] = 32'b11100001100001010111000101000010; //ORR R7 ,R5,R2,ASR #2 //R7 = -123
assign mem[8] = 32'b11100000000001111000000000000011; //AND R8 ,R7,R3 //R8 = -2147483648
assign mem[9] = 32'b11100001111000001001000000000110; //MVN R9 ,R6 //R9 = -11
assign mem[10] = 32'b11100000001001001010000000000101; //EOR R10,R4,R5 //R10 = -84
assign mem[11] = 32'b11100001010110000000000000000110; //CMP R8 ,R6
assign mem[12] = 32'b00010000100000010001000000000001; //ADDNE R1 ,R1,R1 //R1 = 8192
assign mem[13] = 32'b11100001000110010000000000001000; //TST R9 ,R8
assign mem[14] = 32'b00000000100000100010000000000010; //ADDEQ R2 ,R2,R2 //R2 = -1073741824
assign mem[15] = 32'b11100011101000000000101100000001; //MOV R0 ,#1024 //R0 = 1024
assign mem[16] = 32'b11100100100000000001000000000000; //STR R1 ,[R0],#0 //MEM[1024] = 8192
assign mem[17] = 32'b11100100100100001011000000000000; //LDR
assign mem[18] = 32'b11100100100000000010000000000100; //STR R2 ,[R0],#4 //MEM[1028] = -1073741824
assign mem[19] = 32'b11100100100000000011000000001000; //STR R3 ,[R0],#8 //MEM[1032] = -2147483648
assign mem[20] = 32'b11100100100000000100000000001101; //STR R4 ,[R0],#13 //MEM[1036] = 41
assign mem[21] = 32'b11100100100000000101000000010000; //STR R5 ,[R0],#16 //MEM[1040] = -123
assign mem[22] = 32'b11100100100000000110000000010100; //STR R6 ,[R0],#20 //MEM[1044] = 10
assign mem[23] = 32'b11100100100100001010000000000100; //LDR R10,[R0],#4 //R10 = -1073741824
assign mem[24] = 32'b11100100100000000111000000011000; //STR R7 ,[R0],#24 //MEM[1048] = -123
assign mem[25] = 32'b11100011101000000001000000000100; //MOV R1 ,#4 //R1 = 4
assign mem[26] = 32'b11100011101000000010000000000000; //MOV R2 ,#0 //R2 = 0
assign mem[27] = 32'b11100011101000000011000000000000; //MOV R3 ,#0 //R3 = 0
assign mem[28] = 32'b11100000100000000100000100000011; //ADD R4 ,R0,R3,LSL #2
assign mem[29] = 32'b11100100100101000101000000000000; //LDR R5 ,[R4],#0
assign mem[30] = 32'b11100100100101000110000000000100; //LDR R6 ,[R4],#4
assign mem[31] = 32'b11100001010101010000000000000110; //CMP R5 ,R6
assign mem[32] = 32'b11000100100001000110000000000000; //STRGT R6 ,[R4],#0
assign mem[33] = 32'b11000100100001000101000000000100; //STRGT R5 ,[R4],#4
assign mem[34] = 32'b11100010100000110011000000000001; //ADD R3 ,R3,#1
assign mem[35] = 32'b11100011010100110000000000000011; //CMP R3 ,#3
assign mem[36] = 32'b10111010111111111111111111110111; //BLT #-9
assign mem[37] = 32'b11100010100000100010000000000001; //ADD R2 ,R2,#1
assign mem[38] = 32'b11100001010100100000000000000001; //CMP R2 ,R1
assign mem[39] = 32'b10111010111111111111111111110011; //BLT #-13
assign mem[40] = 32'b11100100100100000001000000000000; //LDR R1 ,[R0],#0 //R1 = -2147483648
assign mem[41] = 32'b11100100100100000010000000000100; //LDR R2 ,[R0],#4 //R2 = -1073741824
assign mem[42] = 32'b11100100100100000011000000001000; //LDR R3 ,[R0],#8 //R3 = 41
assign mem[43] = 32'b11100100100100000100000000001100; //LDR R4 ,[R0],#12 //R4 = 8192
assign mem[44] = 32'b11100100100100000101000000010000; //LDR R5 ,[R0],#16 //R5 = -123
assign mem[45] = 32'b11100100100100000110000000010100; //LDR R6 ,[R0],#20 //R4 = 10
assign mem[46] = 32'b11101010111111111111111111111111 ; //B #-


always @(posedge clk, posedge rst) begin
    if(rst) begin
        PC <= 0;
    end
    else if(freeze == 1'b1) begin 
        PC <= PC;
    end
    else begin
        if (Branch_taken == 1'b1)
            PC <= BranchAddr;
        else 
            PC <= PC + 4;
    end
end

assign Instruction = mem[PC >> 2];
endmodule